--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--
--	© 2023 Delta Computer Systems, Inc.
--	Author: Dennis Ritola and David Shroyer
--
--	Additional annotations added by Satchel Hamilton
--
--  Design:         RMC75E Rev 3.n (Replace Xilinx with Microchip)
--  Board:          RMC75E Rev 3.0
--
--	Entity Name		ClockControl
--	File			clockcontrol.vhd
--
--------------------------------------------------------------------------------
--
--	Description: 

	-- The ClockControl module is responsible for controlling the clock signals in the system.
	-- It interfaces with the Clock_Gen component, which generates the clock signals based on the input clock sources.
	-- The module takes various input and output ports, including H1_PRIMARY, H1_CLKWR,
	-- H1_CLK, H1_CLK90, SysClk, RESET, DLL_RST, DLL_LOCK, SysRESET, PowerUp, Enable, and SlowEnable.

	-- Inside the ClockControl module, there are internal signals and processes that handle
	-- the synchronization and control of clock-related operations. These include the synchronization
	-- of the DLL lock status (DLL_LOCK_Int) and the DLL reset command (DLL_RST_sync).
	-- The module also utilizes a one-shot pulse generator (PowerUpOneShot) to generate
	-- initialization pulses on startup or PLL reset. The EnableCount signal is used to
	-- generate enable pulses for clocking the logic at different frequencies.

	-- The module ensures proper synchronization and control of the clock signals
	-- based on the DLL lock status and system reset conditions.
	-- It coordinates the generation and distribution of the
	-- clock signals to different components within the system.

--
--	Revision: 1.3
--
--	File history:
--		Rev 1.3 : 06/08/2023 : 	Added module description
--		Rev 1.2 : 09/01/2022 :	Clean up SysRESET signal
--		Rev 1.1 : 06/10/2022 :	Updated formatting
--
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
-- pragma translate_off
use IEEE.VITAL_Timing.all;
-- pragma translate_on
use IEEE.std_logic_unsigned.all;

-- pragma translate_off
--library unisim;
--use unisim.vcomponents.all;
-- pragma translate_on

entity ClockControl is
	Port ( 
		H1_PRIMARY	: in std_logic;		-- primary clk_in
		H1_CLKWR	: in std_logic;		-- 60MHz input clock for general use
		H1_CLK		: out std_logic;	-- 60MHz system clock 
		H1_CLK90	: out std_logic;	-- 60MHz system clock (90 degree phase lag)
		SysClk		: out std_logic;	-- 30MHz system clock
		RESET		: in std_logic;		-- Sysem reset from power monitor
		DLL_RST		: in std_logic;		-- PLL Reset pulse generated by command from CPU
		DLL_LOCK	: out std_logic;
		SysRESET	: out std_logic;	-- Active when RESET active or PLL not locked
		PowerUp		: out std_logic;
		Enable		: out std_logic;	-- 15.0 MHz system enable (active every 4th 60 MHz clock)
		SlowEnable	: out std_logic		-- 7.5 MHz system enable (active every 8th 60MHz clock)
	);
end ClockControl;

architecture clockcontrol_arch of ClockControl is

	-- Clock_Gen is generated by Microchip's CCC configurator
	component Clock_Gen is
		port (
			-- Inputs
			CLK1_PAD        : in  std_logic;	-- Input 60 MHz clock
			PLL_ARST_N      : in  std_logic;	-- PLL Reset
			PLL_POWERDOWN_N : in  std_logic;	-- PLL Power-down control
			-- Outputs
			GL0             : out std_logic;	-- 60 MHz MDT clock
			GL1             : out std_logic;	-- 60 MHz clock with 90 degree lag
			GL2             : out std_logic;	-- 30 MHz system clock
			LOCK            : out std_logic		-- PLL Locked to within xxx ppm
		);
	end component;

	signal	DLL_LOCK_Int,
			DLLQ1_LOCK		: std_logic;	-- := '0';
	signal	DLL_Lock_ShiftReg	: std_logic_vector (3 downto 0);	-- := x"00000000";
	signal	DLL_Rst_ShiftReg	: std_logic_vector (1 downto 0);	-- := x"00000000";
	signal	DLL_RST_sync	: std_logic;		-- DLL reset command synchronized to system clock
	signal	Reset_int		: std_logic;		-- Flag indicating CPU is ready for FPGA to exit reset
	signal	EnableCount		: std_logic_vector (2 downto 0);	-- := "000";
	signal	PowerUpOneShot	: std_logic_vector (2 downto 0);	-- := "00";
--	signal	sm_cntr			: std_logic_vector (15 downto 0);	-- := x"0000";
--	signal	sm_reset_dcm	: std_logic;	-- := '0';
--	signal	DCM_RESET		: std_logic;	-- := '0';
	
--	signal	TimeCount		: std_logic_vector(25 downto 0);	-- 26 bit counter to generate 1.1 sec delay at 30 MHz
--	signal	DelayDone		: std_logic;						-- Indicates startup delay is done (clock from CPU has had time to change to 60 MHz.)

--	-- State Encoding
--	type STATE_TYPE is array (1 downto 0) of std_logic;
--	constant s0_idle	: STATE_TYPE :="00";
--	constant s1_locked	: STATE_TYPE :="01";
--	constant s2_reset	: STATE_TYPE :="10";
--	constant s3_delay	: STATE_TYPE :="11";
--
--	signal State: STATE_TYPE; -- state can be assigned the constants defined above in "State Encoding"

begin

	-- Note on the commented out sections:
	
	-- This code refers to a previous implementation that is no longer used
	-- in the current design with the Microchip Igloo 2 FPGA.
	
	-- It implements a state machine (StateMachine) that monitors the status of the DLL
	-- (Delay-Locked Loop) and performs certain actions depending on its state.
	-- Here's a breakdown of the commented out code:

	-- The state machine (StateMachine) is a process that is sensitive
	-- to rising edges of the H1_CLKWR signal and the system reset (RESET) signal.

	-- The state machine has four states defined as follows:

	-- s0_idle: Initial state after reset, where the PLL reset signal is kept low.
	-- s1_locked: Monitors the DLL lock status and transitions to the next state if the DLL is not locked.
	-- s2_reset: Resets the DLL for a minimum of three clock cycles.
	-- s3_delay: Waits until the DLL is locked or a delay of 1 millisecond (at 60 MHz) is reached.

	-- Inside the state machine, there are conditions and actions associated with each state:

	-- In the s0_idle state, if the DLL is not locked (DLLQ1_LOCK = '0'), a reset pulse is generated to the DLL.
	-- In the s1_locked state, if the DLL is not locked, a reset pulse is generated to the DLL.
	-- In the s2_reset state, the state machine waits for three clock cycles before transitioning to the s3_delay state.
	-- In the s3_delay state, the state machine waits for either the DLL to lock or a delay of 1 millisecond is reached.
	-- If the delay expires and the DLL is still not locked, it transitions back to the s2_reset state.
	-- If the DLL is locked, it transitions to the s1_locked state.
	
--	-- Monitor PLL for lock. If PLL is not locked, give it a reset signal to attempt to get it to lock.
--	StateMachine : process(H1_CLKWR, RESET)
--	begin
--		if RESET then
--			State <= s0_idle;
--			sm_reset_dcm <= '0';
--		elsif rising_edge(H1_CLKWR) then
--			case State is
--				-- Initial state after reset. Keep PLL reset signal low
--				when s0_idle =>
--					sm_reset_dcm <= '0';
--					-- If PLL is not locked, generate a reset pulse to the PLL
--					if (DLLQ1_LOCK = '0') then
--						sm_cntr(15 downto 0) <= x"0000";
--						sm_reset_dcm <= '1';
--						State <= s2_reset;
--					else
--						State <= s1_locked;
--					end if;
--					
--				-- Monitor for PLL not being locked
--				when s1_locked =>
--					-- If PLL is not locked, generate a reset pulse to the PLL
--					if (DLLQ1_LOCK = '0') then
--						sm_cntr(15 downto 0) <= x"0000";
--						sm_reset_dcm <= '1';
--						State <= s2_reset;
--					end if;
--
--				-- Reset the PLL for a minimum of 3 clock cycles
--				when s2_reset =>
--					if (sm_cntr(15 downto 0) >= x"0004") then
--						sm_cntr(15 downto 0) <= x"0000";
--						sm_reset_dcm <= '0';
--						State <= s3_delay;
--					else
--						sm_cntr(15 downto 0) <= sm_cntr(15 downto 0) + '1';
--					end if;
--
--				-- Wait until PLL locks or for 1 ms.
--				when s3_delay => 
--					if (sm_cntr(15 downto 0) >= x"EA5F") then		-- 1 ms at 60MHz
--						sm_cntr(15 downto 0) <= x"0000";
--						if (DLLQ1_LOCK = '1') then
--							State <= s1_locked;
--						else
--							sm_reset_dcm <= '1';
--							State <= s2_reset;
--						end if;
--					else
--						-- check for lock before delay timer expires
--						if (DLLQ1_LOCK = '1') then
--							sm_cntr(15 downto 0) <= x"0000";
--							State <= s1_locked;
--						else
--							sm_cntr(15 downto 0) <= sm_cntr(15 downto 0) + '1';
--						end if;
--					end if;
--				when others =>	State <= s0_idle;			-- default, reset state
--			end case;
--		end if;
--	end process;

	-- Reset DLL either from a command from CPU or because it is not locked when it should be
--	DCM_RESET <= DLL_RST or sm_reset_dcm;

	-- clkgen was replaced by Microchip's CCC component
	clk_1 : Clock_Gen
		port map (
			-- Inputs
			CLK1_PAD        => H1_PRIMARY,		-- Input 60 MHz clock
--			PLL_ARST_N      => not DCM_RESET,	-- PLL Reset
			PLL_ARST_N      => not RESET,		-- PLL Reset
			PLL_POWERDOWN_N => '1',				-- PLL Power-down control
			-- Outputs
			GL0             => H1_CLK,			-- 60 MHz MDT clock
			GL1             => H1_CLK90,		-- 60 MHz clock with 90 degree lag
			GL2             => SysClk,			-- 30 MHz system clock
			LOCK            => DLLQ1_LOCK		-- PLL Locked to within xxx ppm
		);

	-- The file, discovercontrol.vhd, must also have the FPGA ID byte modified 
	-- to reflect the correct version letter.  ('B' for S/P; 'C' for E)

	-- lock delay shift register
	process (SysClk, RESET)
	begin
		if RESET then
			SysRESET <= '1';
			Reset_int <= '0';
			PowerUpOneShot <= "000";
			PowerUp <= '0';
			DLL_LOCK_Int <= '0';
			DLL_RST_sync <= '0';
			DLL_Lock_ShiftReg <= (others => '0');
			DLL_Rst_ShiftReg <= (others => '0');
			EnableCount <= (others => '0');
			Enable <= '0';
			SlowEnable <= '0';
		elsif rising_edge(SysClk) then
			-- Generate DLL_LOCK signal 4 clock cycles after PLL reports it is locked.
			DLL_Lock_ShiftReg <= DLL_Lock_ShiftReg(2 downto 0) & DLLQ1_LOCK;
			DLL_LOCK_Int <= DLL_Lock_ShiftReg(3) and DLL_Lock_ShiftReg(2) and DLL_Lock_ShiftReg(1) and DLL_Lock_ShiftReg(0);

			-- Synchronize DLL reset command to system clock.
			DLL_Rst_ShiftReg <= DLL_Rst_ShiftReg(0) & DLL_RST;
			DLL_RST_sync <= DLL_Rst_ShiftReg(1);
			
			-- Use the DLL Reset command to set an internal flag indicting CPU is ready for FPGA to come live
			if DLL_RST_sync then
				Reset_int <= '1';
			end if;
			-- If DLL is locked and CPU has commanded a PLL reset then we pull most of the FPGA logic out of reset.
			if Reset_int and DLL_LOCK_Int then
				SysRESET <= '0';
			end if;

			-- Power Up One Shot to generate a single pulse on start-up or PLL reset
			-- This will be used to initialize the control outputs to zero and turn the 
			-- control board LED's to an off state
			PowerUpOneShot <= PowerUpOneShot(1 downto 0) & not SysRESET;
			-- PowerUp pulse generated on rising edge of PowerUpOneShot.
			PowerUp <= not PowerUpOneShot(2) and PowerUpOneShot(1);

			-- Enable Counter to generate an enable pulse every 8th 30MHz clock cycle
			-- this will be used to clock the logic at 7.5MHz and yield a 3.75MHz output clock enable
			-- for the serial data shifting
			EnableCount <= EnableCount + '1';
			if EnableCount(1 downto 0) = "00" then
				Enable <= '1';						-- Active every 133.3ns
			else
				Enable <= '0';
			end if;
			if EnableCount = "000" then
				SlowEnable <= '1';					-- Active every 266.6ns
			else
				SlowEnable <= '0';
			end if;

		end if;
	end process;

	DLL_LOCK <= DLL_LOCK_Int;--LOCKED_delay and DLLQ1_LOCK;

--SysRESET <= RESET or not DLL_LOCK_Int;
--	DLL_LOCK <= DLLQ1_LOCK and DelayDone;--LOCKED_delay and DLLQ1_LOCK;

--	SysRESET <= RESET or not DLLQ1_LOCK or not DelayDone;
--	SysRESET <= RESET or not PowerUpOneShot;
	
--	-- Delay startup until after clock frequency from CPU has been set to 60 MHz. Clock starts off
--	--   at 30 MHz.
--	StartDelay : process (RESET, H1_CLKWR)
--	begin
--		if RESET then
--			TimeCount <= (others => '0');
--			DelayDone <= '0';
--		elsif rising_edge(H1_CLKWR) then
--			if TimeCount(25) = '1' then
--				DelayDone <= '1';
--			else
--				TimeCount <= TimeCount + 1;
--			end if;
--		end if;
--	end process;

end clockcontrol_arch;
