-- Version: 2022.2 2022.2.0.10

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--
--	© 2023 Delta Computer Systems, Inc.
--	Author: SmartDesign
--	
--	Annotations added by Satchel Hamilton
--
--  Design:         RMC75E Rev 3.n (Replace Xilinx with Microchip)
--  Board:          RMC75E Rev 3.0
--
--	Entity Name		Clock_Gen_Clock_Gen_0_FCCC
--	File					Clock_Gen_Clock_Gen_0_FCCC.vhd
--
--------------------------------------------------------------------------------
--
--	Description: 

	-- This module provides the heartbeat of the RMC75E modular motion controller.
	-- It is responsible for generating the raw clock signals used by the rest of the system.
	-- These clock signals are later conditioned to the correct frequencies and phases by the clock_gen module.
	-- The module takes several input and output ports, including LOCK,
	-- PLL_ARST_N, PLL_POWERDOWN_N, CLK1_PAD, and outputs GL0, GL1, and GL2.

	-- Various components are instantiated, such as CLKINT, INBUF, VCC, and GND.
	-- These components handle the buffering, voltage supply, and clock generation functionalities.
	-- The CCC component is also instantiated, which is responsible for generating clock signals with specific configurations.

	-- Overall, the fccc.vhd module forms the initial stage of clock signal generation,
	-- providing the raw clock signals that will be further processed and conditioned in subsequent modules.
	
--	Revision: 1.1
--
--	File history: Rev 1.1 : 06/08/2023 : Added module description
--	
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Clock_Gen_Clock_Gen_0_FCCC is

    port( LOCK            : out   std_logic;
          PLL_ARST_N      : in    std_logic;
          PLL_POWERDOWN_N : in    std_logic;
          CLK1_PAD        : in    std_logic;
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic
        );

end Clock_Gen_Clock_Gen_0_FCCC;

architecture DEF_ARCH of Clock_Gen_Clock_Gen_0_FCCC is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal gnd_net, vcc_net, CLK1_PAD_net, GL0_net, GL1_net, 
        GL2_net : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    GL1_INST : CLKINT
      port map(A => GL1_net, Y => GL1);
    
    CLK1_PAD_INST : INBUF
      port map(PAD => CLK1_PAD, Y => CLK1_PAD_net);
    
    vcc_inst : VCC
      port map(Y => vcc_net);
    
    gnd_inst : GND
      port map(Y => gnd_net);
    
    GL2_INST : CLKINT
      port map(A => GL2_net, Y => GL2);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007DC0000045174001F18C230AC270539DC40404040800101",
         VCOFREQUENCY => 960.000)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => LOCK, BUSY
         => OPEN, CLK0 => vcc_net, CLK1 => vcc_net, CLK2 => 
        vcc_net, CLK3 => vcc_net, NGMUX0_SEL => gnd_net, 
        NGMUX1_SEL => gnd_net, NGMUX2_SEL => gnd_net, NGMUX3_SEL
         => gnd_net, NGMUX0_HOLD_N => vcc_net, NGMUX1_HOLD_N => 
        vcc_net, NGMUX2_HOLD_N => vcc_net, NGMUX3_HOLD_N => 
        vcc_net, NGMUX0_ARST_N => vcc_net, NGMUX1_ARST_N => 
        vcc_net, NGMUX2_ARST_N => vcc_net, NGMUX3_ARST_N => 
        vcc_net, PLL_BYPASS_N => vcc_net, PLL_ARST_N => 
        PLL_ARST_N, PLL_POWERDOWN_N => PLL_POWERDOWN_N, 
        GPD0_ARST_N => vcc_net, GPD1_ARST_N => vcc_net, 
        GPD2_ARST_N => vcc_net, GPD3_ARST_N => vcc_net, PRESET_N
         => gnd_net, PCLK => vcc_net, PSEL => vcc_net, PENABLE
         => vcc_net, PWRITE => vcc_net, PADDR(7) => vcc_net, 
        PADDR(6) => vcc_net, PADDR(5) => vcc_net, PADDR(4) => 
        vcc_net, PADDR(3) => vcc_net, PADDR(2) => vcc_net, 
        PWDATA(7) => vcc_net, PWDATA(6) => vcc_net, PWDATA(5) => 
        vcc_net, PWDATA(4) => vcc_net, PWDATA(3) => vcc_net, 
        PWDATA(2) => vcc_net, PWDATA(1) => vcc_net, PWDATA(0) => 
        vcc_net, CLK0_PAD => gnd_net, CLK1_PAD => CLK1_PAD_net, 
        CLK2_PAD => gnd_net, CLK3_PAD => gnd_net, GL0 => GL0_net, 
        GL1 => GL1_net, GL2 => GL2_net, GL3 => OPEN, 
        RCOSC_25_50MHZ => gnd_net, RCOSC_1MHZ => gnd_net, XTLOSC
         => gnd_net);
end DEF_ARCH; 