--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--
--	© 2023 Delta Computer Systems, Inc.
--	Author: Satchel Hamilton
--
--  Design:         RMC75E Rev 3.n (Replace Xilinx with Microchip)
--  Board:          RMC75E Rev 3.0
--
--	Entity Name		Clock_Gen
--	File			CLK_GEN_NEW.vhd
--
--------------------------------------------------------------------------------
--
--	Description: 
	-- This module generates three clock signals (GL0, GL1, GL2) from an input clock (CLK1_PAD).
	-- The module includes a Phase Locked Loop (PLL) that can be reset (PLL_ARST_N) or powered down (PLL_POWERDOWN_N).
	-- The module also includes a LOCK signal to indicate the status of the PLL.

	-- The primary features of the Clock_Gen module are:
	-- - Generation of a 60MHz clock (GL0) directly derived from the internal clock.
	-- - Generation of a 60MHz clock (GL1) with a 90-degree phase lag relative to GL0. This is achieved using an XOR gate for phase shifting.
	-- - Generation of a 30MHz clock (GL2), which is half the frequency of GL0 and GL1.
	-- - Ability to monitor the status of the PLL via the LOCK signal. The LOCK signal is high when the PLL is neither in reset nor power down mode.

	-- This updated Clock_Gen module replaces two older modules that were affected by a compatibility issue between ModelSim and SmartFusion2.
	-- The issues related to the compatibility have been addressed in this module.
	-- However, the new module maintains the same interface and functionality, providing a drop-in replacement for the older modules.

	-- Ports:
	-- - Inputs:
	  -- - CLK1_PAD: The primary external clock input.
	  -- - PLL_ARST_N: System reset from power monitor.
	  -- - PLL_POWERDOWN_N: PLL Reset pulse generated by command from CPU.
	-- - Outputs:
	  -- - GL0: 60MHz system clock.
	  -- - GL1: 60MHz system clock with 90 degree phase lag.
	  -- - GL2: 30MHz system clock.
	  -- - LOCK: PLL lock signal.

	-- Reset and Power Down:
	-- - If PLL_ARST_N is high, or if PLL_POWERDOWN_N is high, the internal clock is reset.
	-- - The LOCK signal is high when the PLL is neither in reset nor in power down mode.

	-- Architecture:
	-- - The architecture of this module (Behavioral) implements clock signal generation using a series
	-- of processes that trigger on either the rising edge of the external or internal clocks.

	-- Compatibility:
	-- - This module has been tested for compatibility with the ModelSim environment and RMC75E source code.

	-- Note: For the accurate simulation of the module, the external CLK1_PAD signal should be a 120MHz clock
	-- for the generated clocks to have the specified frequencies.

--	Revision: 1.0
--
--	File history:
--	
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity Clock_Gen is
    port( 
        CLK1_PAD           : in  std_logic;  -- primary clk_in
        PLL_ARST_N         : in  std_logic;  -- System reset from power monitor
        PLL_POWERDOWN_N    : in  std_logic;  -- PLL Reset pulse generated by command from CPU
        -- Outputs
        GL0                : out std_logic;  -- 60MHz system clock 
        GL1                : out std_logic;  -- 60MHz system clock (90 degree phase lag)
        GL2                : out std_logic;  -- 30MHz system clock
        LOCK               : out std_logic   -- PLL lock signal
    );
end Clock_Gen;

architecture Behavioral of Clock_Gen is
    signal internal_clock: std_logic;
    signal phase_shift_clock: std_logic;
    signal clk_60MHz: std_logic := '0';
    signal clk_60MHz_90deg: std_logic := '0';
    signal clk_30MHz: std_logic := '0';

begin
    -- main clock process
    clock_process : process(CLK1_PAD)
    begin
        if rising_edge(CLK1_PAD) then
            if PLL_ARST_N = '1' then
                internal_clock <= '0';
            elsif PLL_POWERDOWN_N = '1' then
                internal_clock <= '0';
            else
                internal_clock <= not internal_clock;
            end if;
        end if;
    end process clock_process;

    -- generate 60MHz clock
    clk_60MHz_gen : process(internal_clock)
    begin
        if rising_edge(internal_clock) then
            clk_60MHz <= not clk_60MHz;
        end if;
    end process clk_60MHz_gen;

    -- generate 60MHz clock with 90 degree phase shift using XOR gate
    clk_60MHz_90deg_gen : process(internal_clock, clk_60MHz)
    begin
        clk_60MHz_90deg <= internal_clock xor clk_60MHz;
    end process clk_60MHz_90deg_gen;

    -- generate 30MHz clock
    clk_30MHz_gen : process(clk_60MHz)
    begin
        if rising_edge(clk_60MHz) then
            clk_30MHz <= not clk_30MHz;
        end if;
    end process clk_30MHz_gen;

    -- output signals
    GL0 <= clk_60MHz;
    GL1 <= clk_60MHz_90deg;
    GL2 <= clk_30MHz;
    LOCK <= not PLL_ARST_N and not PLL_POWERDOWN_N;  -- simplified, indicates it's not in reset or powerdown
end Behavioral;
