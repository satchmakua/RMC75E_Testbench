--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--
--	© 2022 Delta Computer Systems, Inc.
--	Author: Dennis Ritola and David Shroyer
--
--	Design:			RMC75E Rev 3.n (Replace Xilinx with Microchip)
--	Board:			RMC75E Rev 3.0
--
--	Entity Name		CPUConfig
--	File			CPUConfig.vhd
--
--------------------------------------------------------------------------------
--
--	Description: 
--		
--
--	Revision: 1.1
--
--	File history:
--		Rev 1.1 : 06/07/2022 :	Updated formatting
--
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CPUConfig is
	Port (
		RESET				: in std_logic;		-- External Reset from power monitor and watchdog IC.
		SysRESET			: in std_logic;		-- Main internal reset. Used to clear DLL_RST
		H1_CLKWR			: in std_logic;
		H1_PRIMARY			: in std_logic;							-- 60MHz system clock
		intDATA				: in std_logic_vector (31 downto 0);
		cpuConfigDataOut	: out std_logic_vector (31 downto 0);
		CPUConfigWrite		: in std_logic;
		M_DRV_EN_L			: out std_logic;						-- Control Output Enable Line
		HALT_DRIVE_L		: in std_logic;
		DLL_LOCK			: in std_logic;
		DLL_RST				: out std_logic;	-- Was for resetting DLL. Now used to clear SysRESET. Generated by command from CPU.
		LoopTime			: out std_logic_vector (2 downto 0);	-- Control Loop Time Selection
		ENET_Build			: in std_logic
	);
end CPUConfig;

architecture CPUConfig_arch of CPUConfig is

	signal	int_M_DRV_EN,
			int_DLL_RST			: std_logic;	-- := '0';
	signal	intLoopTime			: std_logic_vector (2 downto 0);	-- := "000";
	signal	dll_rst_pre_queue	: std_logic;	-- := '0';
	signal	dll_rst_queue		: std_logic_vector (1 downto 0);	-- := x"00";

begin

	LoopTime(2 downto 0) <= intLoopTime(2 downto 0);

	cpuConfigDataOut(31 downto 0) <= "0000000000000000000000000" & intLoopTime(2 downto 0) & '0' & '0' & DLL_LOCK & int_M_DRV_EN;

	-- The actual drive enable line is active low. The power-up default 
	-- condition is off. The processor will write to the bit as if it's 
	-- active high. 
	process (RESET, H1_CLKWR)
	begin
		if RESET then
			int_M_DRV_EN <= '0';    -- whenever a power dip/drop is detected, kill the drives
		elsif rising_edge(H1_CLKWR) then
			if HALT_DRIVE_L = '0' then
				int_M_DRV_EN <= '0';    -- whenever a power dip/drop is detected, kill the drives
			elsif CPUConfigWrite = '1' then
				int_M_DRV_EN <= intDATA(0);
			end if;

			if CPUConfigWrite = '1' then
--				PROFIEnable <= intDATA(3) and not ENET_Build;
				intLoopTime(2 downto 0) <= intDATA(6 downto 4);
			end if;
		end if;
	end process;

	M_DRV_EN_L <= not int_M_DRV_EN;

	process (RESET, H1_PRIMARY)
	begin
		if RESET then
			int_DLL_RST <= '0';
			DLL_RST <= '0';
			dll_rst_pre_queue <= '0';
			dll_rst_queue <= (others => '0');
		elsif rising_edge(H1_PRIMARY) then
			-- Once the SysRESET is low, clear DLL_RST (which is the signal used to set SysRESET low)
			if not SysRESET then
				int_DLL_RST <= '0';
			-- If SysRESET is high, a write to bit 2 will generate a DLL_RST signal used now to clear internal reset (SysRESET)
			elsif CPUConfigWrite = '1' then
				int_DLL_RST <= intDATA(2);
			end if;

			-- This added level of protection ensures that no glitches sneak through during the write process
			-- The DLL reset is quite sensitive to these small glitches and the effect is catastrophic to the FPGA.
			if CPUConfigWrite = '0' then
				dll_rst_pre_queue <= int_DLL_RST;
			end if;

			dll_rst_queue(1 downto 0) <= dll_rst_queue(0) & dll_rst_pre_queue;

			DLL_RST <= dll_rst_queue(1);

		end if;
	end process;

end CPUConfig_arch;
